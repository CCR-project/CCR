Require Import Coqlib.
Require Import ITreelib.
Require Import Universe.
Require Import Skeleton.
Require Import PCM.

Set Implicit Arguments.


Section EVENTS.

  Inductive eventE: Type -> Type :=
  | Choose X: eventE X
  | Take X: eventE X
  | Syscall (fn: fname) (m: Mem.t) (args: list val): eventE (Mem.t * val)
  (*** Syscall should be able to look at current memory (full information).
       Normal modules will call Memory (Language) module in order to call system call,
       because Memory (Language) module is the only one with access to Mem.t.
   ***)
  .

  Inductive callE: Type -> Type :=
  | Call (fn: fname) (args: list val): callE val
  .

  (* Notation "'Choose' X" := (trigger (Choose X)) (at level 50, only parsing). *)
  (* Notation "'Take' X" := (trigger (Take X)) (at level 50, only parsing). *)

  Definition triggerUB {E A} `{eventE -< E}: itree E A :=
    v <- trigger (Take void);; match v: void with end
  .

  Definition triggerNB {E A} `{eventE -< E}: itree E A :=
    v <- trigger (Choose void);; match v: void with end
  .

  Definition unwrapN {E X} `{eventE -< E} (x: option X): itree E X :=
    match x with
    | Some x => ret x
    | None => triggerNB
    end.

  Definition unwrapU {E X} `{eventE -< E} (x: option X): itree E X :=
    match x with
    | Some x => ret x
    | None => triggerUB
    end.

  Definition assume {E} `{eventE -< E} (P: Prop): itree E unit := trigger (Take P) ;; Ret tt.
  Definition guarantee {E} `{eventE -< E} (P: Prop): itree E unit := trigger (Choose P) ;; Ret tt.

  (* Notation "'unint?'" := (unwrapA <*> unint) (at level 57, only parsing). *)
  (* Notation "'unint﹗'" := (unwrapG <*> unint) (at level 57, only parsing). *)
  (* Notation "'Ret!' f" := (RetG f) (at level 57, only parsing). *)
  (* Notation "'Ret?' f" := (RetA f) (at level 57, only parsing). *)

  Context `{GRA: GRA.t}.

  Inductive rE: Type -> Type :=
  (* | MPut (mn: mname) (r: GRA): rE unit *)
  (* | MGet (mn: mname): rE GRA *)
  (* | FPut (r: GRA): rE unit *)
  (* | FGet: rE GRA *)
  | Put (mn: mname) (mr: GRA) (fr: GRA): rE unit
  | MGet (mn: mname): rE GRA
  | FGet: rE GRA
  (* | Get (mn: mname): rE (GRA * GRA) *)

  (*** NOTE: These methods can be implemented using Put/Get,
       but making it explicit will be helpful for meta-theory.
       E.g., In top-level, if all modules are well-typed,
       we can make "CheckWf" to Nop by adjusting handler.
   ***)
  | Forge (fr: GRA): rE unit
  | Discard (fr: GRA): rE unit
  | CheckWf (mn: mname): rE unit

  | PushFrame: rE unit
  | PopFrame: rE unit
  .

  Definition MPut E `{rE -< E} (mn: mname) (mr: GRA): itree E unit :=
    fr <- trigger FGet;;
    trigger (Put mn mr fr)
  .

  (*** TODO: we don't want to require "mname" here ***)
  (*** use dummy mname? ***)
  (* Definition FPut E `{rE -< E} (mn: mname) (fr: GRA): itree E unit := *)

  Definition Es: Type -> Type := (callE +' rE +' eventE).

  (* Inductive mdE: Type -> Type := *)
  (* | MPut (mn: mname) (r: GRA): mdE unit *)
  (* | MGet (mn: mname): mdE GRA *)
  (* . *)

  (* Inductive fnE: Type -> Type := *)
  (* | FPut (r: GRA): fnE unit *)
  (* | FGet: fnE GRA *)
  (* | FPush: fnE unit *)
  (* | FPop: fnE unit *)
  (* . *)

End EVENTS.

Notation "f '?'" := (unwrapU f) (at level 60, only parsing).
Notation "f '﹗'" := (unwrapN f) (at level 60, only parsing).





Module ModSem.
Section MODSEM.

  (* Record t: Type := mk { *)
  (*   state: Type; *)
  (*   local_data: Type; *)
  (*   step (skenv: SkEnv.t) (st0: state) (ev: option event) (st1: state): Prop; *)
  (*   state_sort: state -> sort; *)
  (*   initial_local_data: local_data; *)
  (*   sk: Sk.t; *)
  (*   name: string; *)
  (* } *)
  (* . *)

  Context `{GRA: GRA.t}.

  Record t: Type := mk {
    sk: Sk.t;
    (* initial_ld: mname -> GRA; *)
    sem: callE ~> itree Es;
    initial_ld: list (mname * GRA);
  }
  .

  Definition wf (md: t): Prop := Sk.wf md.(sk).

  (*** using "Program Definition" makes the definition uncompilable; why?? ***)
  Definition merge (md0 md1: t): t := {|
    sk := Sk.add md0.(sk) md1.(sk);
    (* initial_ld := URA.add (t:=URA.pointwise _ _) md0.(initial_ld) md1.(initial_ld); *)
    sem := fun _ '(Call fn args) =>
             (if List.in_dec string_dec fn md0.(sk) then md0.(sem) else md1.(sem)) _ (Call fn args);
    initial_ld := app md0.(initial_ld) md0.(initial_ld);
  |}
  .

End MODSEM.
End ModSem.



Inductive pred: Type :=
| true
| false
| meta (P: Prop)

| disj: pred -> pred -> pred
| conj: pred -> pred -> pred
| neg: pred -> pred
| impl: pred -> pred -> pred

| univ (X: Type): (X -> pred) -> pred
| exst (X: Type): (X -> pred) -> pred
.

(*** https://en.wikipedia.org/wiki/Negation_normal_form ***)
Fixpoint embed (p: pred): itree eventE unit :=
  match p with
  | true => triggerUB
  | false => triggerNB
  | meta P => guarantee P

  | disj p0 p1 => b <- trigger (Choose _);; if (b: bool) then embed p0 else embed p1
  | conj p0 p1 => b <- trigger (Take _);; if (b: bool) then embed p0 else embed p1
  | neg p =>
    match p with
    | meta P => assume P
    | _ => triggerNB (*** we are assuming negation normal form ***)
    end
  | impl _ _ => triggerNB (*** we are assuming negation normal form ***)

  | @univ X k => x <- trigger (Take X);; embed (k x)
  | @exst X k => x <- trigger (Choose X);; embed (k x)
  end
.

(*** TODO: implication --> function call? ***)
(***
P -> Q
~=
pname :=
  embed P

pqname :=
  (call pname) (finite times);;
  embed Q




(P -> Q) -> R
~=
pname :=
  embed P

pqname :=
  (call pname) (finite times);;
  embed Q

pqrname :=
  (call pqname) (finite times);;
  embed R
***)

(* Fixpoint embed (p: pred) (is_pos: bool): itree eventE unit := *)
(*   match p with *)
(*   | true => triggerUB *)
(*   | false => triggerNB *)
(*   | meta P => guarantee P *)
(*   | disj p0 p1 => b <- trigger (Choose _);; if (b: bool) then embed p0 is_pos else embed p1 is_pos *)
(*   | conj p0 p1 => b <- trigger (Take _);; if (b: bool) then embed p0 is_pos else embed p1 is_pos *)
(*   | @univ X k => x <- trigger (Take X);; embed (k x) is_pos *)
(*   | @exst X k => x <- trigger (Choose X);; embed (k x) is_pos *)
(*   | _ => triggerNB *)
(*   end *)
(* . *)
